lpm_mux20_inst : lpm_mux20 PORT MAP (
		data0x	 => data0x_sig,
		data1x	 => data1x_sig,
		data2x	 => data2x_sig,
		sel	 => sel_sig,
		result	 => result_sig
	);
